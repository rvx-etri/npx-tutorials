`ifndef __DCA_MATRIX_INFO_H__
`define __DCA_MATRIX_INFO_H__

`include "dca_matrix_info_memorymap_offset.vh"

`define GEN_DCA_DCA_MATRIX_DATATYPE(is_float, is_signed, addr_lsa, num_bits) (((addr_lsa&0x07)<<2)|((is_float&0x1)<<1)|((is_signed&0x1)<<0))

`define DCA_MATRIX_DATATYPE_UINT01 GEN_DCA_MATRIX_DATATYPE(0,0,-3,1)
`define DCA_MATRIX_DATATYPE_SINT02 GEN_DCA_MATRIX_DATATYPE(0,1,-2,2)
`define DCA_MATRIX_DATATYPE_UINT02 GEN_DCA_MATRIX_DATATYPE(0,0,-2,2)
`define DCA_MATRIX_DATATYPE_SINT04 GEN_DCA_MATRIX_DATATYPE(0,1,-1,4)
`define DCA_MATRIX_DATATYPE_UINT04 GEN_DCA_MATRIX_DATATYPE(0,0,-1,4)
`define DCA_MATRIX_DATATYPE_SINT08 GEN_DCA_MATRIX_DATATYPE(0,1,0,8)
`define DCA_MATRIX_DATATYPE_UINT08 GEN_DCA_MATRIX_DATATYPE(0,0,0,8)
`define DCA_MATRIX_DATATYPE_SINT16 GEN_DCA_MATRIX_DATATYPE(0,1,1,16)
`define DCA_MATRIX_DATATYPE_UINT16 GEN_DCA_MATRIX_DATATYPE(0,0,1,16)
`define DCA_MATRIX_DATATYPE_SINT32 GEN_DCA_MATRIX_DATATYPE(0,1,2,32)
`define DCA_MATRIX_DATATYPE_FLOAT32 GEN_DCA_MATRIX_DATATYPE(1,1,2,32)

`define BW_DCA_MATRIX_INFO (`BW_DCA_MATRIX_INFO_ADDR+`BW_DCA_MATRIX_INFO_STRIDE_LS3+`BW_DCA_MATRIX_INFO_NUM_ROW_M1+`BW_DCA_MATRIX_INFO_NUM_COL_M1+`BW_DCA_MATRIX_INFO_IS_SIGNED+`BW_DCA_MATRIX_INFO_IS_FLOAT+`BW_DCA_MATRIX_INFO_ADDR_LSA_P3)

`define BW_DCA_MATRIX_INFO_ALIGNED ((((`BW_DCA_MATRIX_INFO-1)>>5)+1)<<5)

`endif
